module counter(out, clk, reset);
	parameter WIDTH = 8;
	output [WIDTH-1 : 0] out;
	input clk, reset;
endmodule
